/* Package: rvt_pkg
 * Includes all RiVET base objects.
 */
package rvt_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "dv_macros.svh"
  `include "rvt_macros.svh"

  typedef enum int {
    SubNone,
    SubChecker,
    SubCoverage,
    SubLogger
  } sub_mode_e;

  `include "rvt_base_obj.svh"
  `include "rvt_base_cmp.svh"

  `include "rvt_base_item.svh"
  `include "rvt_base_agnt.svh"

  `include "rvt_bfm_cb.svh"
  `include "rvt_bfm.svh"

  `include "rvt_core_cfg.svh"

  `include "rvt_cfg.svh"
  `include "rvt_agent_cfg.svh"

  `include "rvt_seqr.svh"

  `include "rvt_sequence.svh"

  `include "rvt_monitor.svh"
  `include "rvt_driver.svh"
  `include "rvt_subscriber.svh"

  `include "rvt_base_agent.svh"
  `include "rvt_agent.svh"
endpackage : rvt_pkg
