package tev_verif_pkg;


    // Base Items
    `include "tev_base_config_c.svh"
    `include "tev_base_tem_c.svh"
    `include "tev_base_compnent_c.svh"
endpackage
