/**
 * @class rvt_instr
 * RISC-V instruction object.
 * Contains all coverage and randomization related utilities.
 */

`ifndef _RVT_INSTR_
`define _RVT_INSTR_
class rvt_instr_cov extends rvt_obj;

endclass : rvt_instr_cov
`endif //_RVT_INSTR_
