package rvt_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "dv_macros.svh"

  import rvt_base_pkg::*;
  import rvt_mem_pkg::*;
endpackage
