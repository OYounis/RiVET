package rvt_mem_pkg;
  import uvm_pkg::*;
  import rvt_base_pkg::*;
  `include"uvm_macros.svh"

  `include "rvt_mem_cfg.svh"
  `include "rvt_mem_item.svh"
  `include "rvt_mem.svh"
  `include "rvt_mem_sequencer.svh"
  `include "rvt_mem_driver.svh"
  `include "rvt_mem_monitor.svh"
  `include "rvt_mem_agent.svh"

  `include "rvt_mem_sequence.svh"
endpackage : rvt_mem_pkg
