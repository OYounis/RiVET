class tev_base_item_c extends uvm_sequence_item;
    `uvm_object_utils(tev_base_item_c)

    function new(string name = "tev_base_item");
        super.new(name);
    endfunction

endclass
