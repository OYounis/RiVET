
package rvt_core_pkg;
endpackage : rvt_core_pkg
