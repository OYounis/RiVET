class tev_instr_item_c extends tev_base_item_c;
    `uvm_object_utils(tev_instr_item_c)
    function new(string name = "tev_instr_item");
        super.new(name);
    endfunction
endclass
